/******************************************************************************
 *     "Copyright (C) 2014, Codasip s.r.o., All Rights Reserved"              *
 ******************************************************************************/
/**
 *  \file
 *  \date   Sat Jul 19 17:47:35 2014
 *  \author Codasip HW generator v2.2.0.internal
 *  \brief  Definition of the 'sv_codix_risc_platform_ca_t_gm_pkg' package.
 */

package sv_codix_risc_platform_ca_t_gm_pkg;
	import uvm_pkg::*;
	import sv_param_pkg::*;
	import sv_codix_risc_ca_t_agent_pkg::*;
	import sv_codix_risc_platform_ca_t_agent_pkg::*;
	import codix_risc_platform_ia_dpi_pkg::*;

	`include "uvm_macros.svh"
	`include "golden_model.svh"
endpackage: sv_codix_risc_platform_ca_t_gm_pkg
