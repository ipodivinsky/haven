--  ---------------------------------------------------------
--  Hardware Accelerated Functional Verification of Processor
--  ---------------------------------------------------------

--  \file   program_driver.vhd
--  \date   29-04-2014
--  \brief  Testbench for testing program driver
--  \author Jakub Podivinsky, ipodivinsky@fit.vutbr.cz
--
--  \input  Input signals for program driver are generated by 
--          FL_BFM component by function: 
--          SendWriteFile("path to input data file", EVER, flCmd_0, 0);
--
--          Format of "input data file" is following: 
--             00000000 --start header
--             00000001
--             #
--             00000000 --data header
--             00000000
--             instruction 0
--             instruction 1
--             instruction 2
--                   .
--                   .
--                   .
--             instruction n
--             # 
--             00000000 --data header
--             00000000 --it is posibble to send new data packet before stop header
--             instruction n+1 --also it is available to send new data packet before stop header from other file
--             instruction n+2
--                   .
--                   .
--                   .
--             instruction n +m
--             #
--             00000000 --stop header
--             00000004 --after stop header it is imposibble to send new data packet
--             #
--
--          Example of input file:
--             ./input/test_simple - simple set of instructions
--             ./input/test_1half - simple set of instructions without stop header
--             ./input/test_2half - simple set of instruction without start header
--             ./input/full_program - real program
--

library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.fl_sim_oper.all;
use work.fl_bfm_pkg.all;
use work.fl_bfm_rdy_pkg.all;


entity testbench is
end entity testbench;

architecture behavioral of testbench is

   -- constants
   constant IN_DATA_WIDTH        : integer := 64;
   constant OUT_DATA_WIDTH       : integer := 32;

   constant clkper               : time := 10 ns; 
   constant reset_time           : time := 100 ns;

   -- signals
   signal clk                    : std_logic;
   signal reset                  : std_logic;
   
   -- UUT input signals
   signal driver_in_data         : std_logic_vector(IN_DATA_WIDTH-1 downto 0);
   signal driver_in_rem          : std_logic_vector(2 downto 0);
   signal driver_in_sof_n        : std_logic;
   signal driver_in_sop_n        : std_logic;
   signal driver_in_eof_n        : std_logic;
   signal driver_in_eop_n        : std_logic;
   signal driver_in_src_rdy_n    : std_logic;
   signal driver_in_dst_rdy_n    : std_logic;
   signal driver_in_mem_done     : std_logic;
   
   -- UUT output signals
   signal driver_out_done        : std_logic;
   signal driver_proc_reset      : std_logic;
   signal driver_out_d0          : std_logic_vector(OUT_DATA_WIDTH-1 downto 0);
   signal driver_out_dbg_mode    : std_logic;
   signal driver_out_wa0         : std_logic_vector(18 downto 0);
   signal driver_out_we0         : std_logic;
   signal driver_out_wsc0        : std_logic_vector(2 downto 0);
   signal driver_out_wsi0        : std_logic_vector(1 downto 0);

-- ----------------------------------------------------------------------------
--                      Architecture body
-- ----------------------------------------------------------------------------
begin

   -- -------------------------------------------------------------------------
   --                   program driver
   -- -------------------------------------------------------------------------
   uut: entity work.PROGRAM_DRIVER
      generic map (
         IN_DATA_WIDTH     => IN_DATA_WIDTH,
         OUT_DATA_WIDTH    => OUT_DATA_WIDTH
      )
      port map (
         CLK               => clk,
         RESET             => reset,

         RX_DATA           => driver_in_data,
         RX_REM            => driver_in_rem,
         RX_SOF_N          => driver_in_sof_n,
         RX_SOP_N          => driver_in_sop_n,
         RX_EOP_N          => driver_in_eop_n,
         RX_EOF_N          => driver_in_eof_n,
         RX_SRC_RDY_N      => driver_in_src_rdy_n,
         RX_DST_RDY_N      => driver_in_dst_rdy_n,

         MEM_DONE          => driver_in_mem_done,
         DONE              => driver_out_done,
         
         proc_reset        => driver_proc_reset,
         
         dbg_mode_mem_D0   => driver_out_d0,
         dbg_mode_mem      => driver_out_dbg_mode,
         dbg_mode_mem_WA0  => driver_out_wa0,
         dbg_mode_mem_WE0  => driver_out_we0,
         dbg_mode_mem_WSC0 => driver_out_wsc0,
         dbg_mode_mem_WSI0 => driver_out_wsi0

      );
	  
   -- -------------------------------------------------------------------------
   --                           Input FL_BFM
   -- -------------------------------------------------------------------------
   FL_BFM_I: entity work.FL_BFM
   generic map (
      DATA_WIDTH => IN_DATA_WIDTH,
      FL_BFM_ID => 00
   )
   port map (
      -- Common interface
      RESET           => reset,
      CLK             => clk,

      TX_DATA         => driver_in_data,
      TX_REM          => driver_in_rem,
      TX_SOF_N        => driver_in_sof_n,
      TX_EOF_N        => driver_in_eof_n,
      TX_SOP_N        => driver_in_sop_n,
      TX_EOP_N        => driver_in_eop_n,
      TX_SRC_RDY_N    => driver_in_src_rdy_n,
      TX_DST_RDY_N    => driver_in_dst_rdy_n
   ); 
   
   -- -------------------------------------------------------------------------
   --                           CLK generator
   -- -------------------------------------------------------------------------
   clkgen: process
   begin
      clk <= '1';
      wait for clkper/2;
      clk <= '0';
      wait for clkper/2;
   end process;

   -- -------------------------------------------------------------------------
   --                           RESET generator
   -- -------------------------------------------------------------------------   
   resetgen: process
   begin
      reset <= '1';
      wait for reset_time;
      reset <= '0';
      wait;
   end process;

   -- -------------------------------------------------------------------------
   --                           Testbech process
   -- -------------------------------------------------------------------------   
   tb: process

   begin

      driver_in_mem_done <= '0';
      wait for reset_time; 
      wait until rising_edge(clk);
      
      SendWriteFile("./input/test_1half", EVER, flCmd_0, 0);
      --SendWriteFile("./input/test_simple", EVER, flCmd_0, 0);
      --SendWriteFile("./input/full_program", EVER, flCmd_0, 0);
      
	  
      wait until rising_edge(clk);
      
      SendWriteFile("./input/test_2half", EVER, flCmd_0, 0);
      
      wait until rising_edge(clk);
      wait until rising_edge(clk);
      wait until rising_edge(clk);
     
      driver_in_mem_done <= '1'; 
	  
      wait until rising_edge(clk);
      wait until rising_edge(clk);
      
      driver_in_mem_done <= '0';
	  
      
      SendWriteFile("./input/test_simple", EVER, flCmd_0, 0);
      wait;
      
  end process tb; 
   
end architecture behavioral;
