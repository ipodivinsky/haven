/******************************************************************************
 *     "Copyright (C) 2014, Codasip s.r.o., All Rights Reserved"              *
 ******************************************************************************/
/**
 *  \file
 *  \date   Sat Jul 19 17:47:35 2014
 *  \author Codasip HW generator v2.2.0.internal
 *  \brief  Definition of the 'sv_codix_risc_ca_core_main_instr_hw_instr_hw_t_agent_pkg' package.
 */

package sv_codix_risc_ca_core_main_instr_hw_instr_hw_t_agent_pkg;
	import uvm_pkg::*;
	import sv_param_pkg::*;

	`include "uvm_macros.svh"
	`include "decoder.svh"
	`include "transaction.svh"
	`include "ifc_wrapper.svh"
	`include "config.svh"
	`include "monitor.svh"
	`include "coverage.svh"
	`include "agent.svh"
endpackage: sv_codix_risc_ca_core_main_instr_hw_instr_hw_t_agent_pkg
