--  ---------------------------------------------------------
--  Hardware Accelerated Functional Verification of Processor
--  ---------------------------------------------------------

--  \file   program_driver.vhd
--  \date   05-05-2014
--  \brief  Testbench for testing verification core
--  \author Jakub Podivinsky, ipodivinsky@fit.vutbr.cz
--
--  \input  Input signals for verification core are generated by 
--          FL_BFM component by function: 
--          SendWriteFile("path to input data file", EVER, flCmd_0, 0);
--
--          Format of "input data file" is following: 
--             00000000 --start header
--             00000001
--             #
--             00000000 --data header
--             00000000
--             instruction 0
--             instruction 1
--             instruction 2
--                   .
--                   .
--                   .
--             instruction n
--             # 
--             00000000 --data header
--             00000000 --it is posibble to send new data packet before stop header
--             instruction n+1 --also it is available to send new data packet before stop header from other file
--             instruction n+2
--                   .
--                   .
--                   .
--             instruction n +m
--             #
--             00000000 --stop header
--             00000004 --after stop header it is imposibble to send new data packet
--             #
--
--          Example of input file:
--             ./input/input_program_hex - real program
--
--  \output Output FrameLink protocol signals are processed by 
--          FL_MONITOR component, data are store in file ./output/monitor 
--
--          Format of output file: 
--             00000001    -- header [7..0]
--             00000000    -- header [15..8]
--             .DATA 0.    -- data [7..0]
--             #           -- end of packet
--             00000001    
--             00000000    
--             .DATA 1.   
--             #    
--                .
--                .
--                .
--             00000001    
--             00000000    
--             .DATA n.   
--             #   

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use work.fl_sim_oper.all;
use work.fl_bfm_pkg.all;
use work.fl_bfm_rdy_pkg.all;

library work;

-- HAVEN constants
use work.haven_const.all;

entity testbench is
end entity;

architecture test of testbench is

   -- ------------------------------------------------------------------------
   --                                Constants
   -- ------------------------------------------------------------------------

   -- data width
   constant FL_DATA_WIDTH      : integer := 64; -- FrameLink data width
   constant CODIX_DATA_WIDTH   : integer := 32; -- processor data width

   -- duration of reset
   constant RESET_TIME  : time := 100 ns;
   -- clock period
   constant CLK_PERIOD  : time := 10 ns;

   -- ------------------------------------------------------------------------
   --                                 Signals
   -- ------------------------------------------------------------------------

   -- common signals
   signal clk           : std_logic;
   signal reset         : std_logic;

   -- input FrameLink
   signal rx_data       : std_logic_vector(FL_DATA_WIDTH-1 downto 0);
   signal rx_rem        : std_logic_vector(2 downto 0);
   signal rx_sof_n      : std_logic;
   signal rx_eof_n      : std_logic;
   signal rx_sop_n      : std_logic;
   signal rx_eop_n      : std_logic;
   signal rx_src_rdy_n  : std_logic;
   signal rx_dst_rdy_n  : std_logic;

   -- output FrameLink
   signal tx_data       : std_logic_vector(FL_DATA_WIDTH-1 downto 0);
   signal tx_rem        : std_logic_vector(2 downto 0);
   signal tx_sof_n      : std_logic;
   signal tx_eof_n      : std_logic;
   signal tx_sop_n      : std_logic;
   signal tx_eop_n      : std_logic;
   signal tx_src_rdy_n  : std_logic;
   signal tx_dst_rdy_n  : std_logic;

   -- MI32 interface
   signal mi32_dwr      : std_logic_vector(31 downto 0);
   signal mi32_addr     : std_logic_vector(31 downto 0);
   signal mi32_rd       : std_logic;
   signal mi32_wr       : std_logic;
   signal mi32_be       : std_logic_vector(3 downto 0);
   signal mi32_drd      : std_logic_vector(31 downto 0);
   signal mi32_ardy     : std_logic;
   signal mi32_drdy     : std_logic;

--   -- Reverse function to change bit-order inside byte.
--   function reverse( src: std_logic_vector ) return std_logic_vector is
--      variable result: std_logic_vector( src'range );
--      alias r_src: std_logic_vector( src'reverse_range ) is src;
--      begin
--         for ii in r_src'range loop
--            result(ii) := r_src(ii);
--         end loop;
--         return result;
--   end function;

begin

   -- -----------------------------------------------------------------------
   --                             Unit under test
   -- -----------------------------------------------------------------------
   uut: entity work.verification_core
   generic map(
      -- data width 
      FL_DATA_WIDTH      => FL_DATA_WIDTH, -- FrameLink data width
      CODIX_DATA_WIDTH   => CODIX_DATA_WIDTH, -- processor data width
      -- the CORE_TYPE generic specifies the verified unit in the core
      CORE_TYPE          => codasip_codix
   )
   port map(
      CLK            => clk,
      RESET          => reset,

      -- FrameLink input interface
      RX_DATA        => rx_data,
      RX_REM         => rx_rem,
      RX_SOF_N       => rx_sof_n,
      RX_EOF_N       => rx_eof_n,
      RX_SOP_N       => rx_sop_n,
      RX_EOP_N       => rx_eop_n,
      RX_SRC_RDY_N   => rx_src_rdy_n,
      RX_DST_RDY_N   => rx_dst_rdy_n,

      -- FrameLink output interface
      TX_DATA        => tx_data,
      TX_REM         => tx_rem,
      TX_SOF_N       => tx_sof_n,
      TX_EOF_N       => tx_eof_n,
      TX_SOP_N       => tx_sop_n,
      TX_EOP_N       => tx_eop_n,
      TX_SRC_RDY_N   => tx_src_rdy_n,
      TX_DST_RDY_N   => tx_dst_rdy_n,

      -- MI32 interface (actually unused)
      MI32_DWR       => mi32_dwr,
      MI32_ADDR      => mi32_addr,
      MI32_RD        => mi32_rd,
      MI32_WR        => mi32_wr,
      MI32_BE        => mi32_be,
      MI32_DRD       => mi32_drd,
      MI32_ARDY      => mi32_ardy,
      MI32_DRDY      => mi32_drdy

   );

   -- -------------------------------------------------------------------------
   --                           Input FL_BFM
   -- -------------------------------------------------------------------------
   FL_BFM_I: entity work.FL_BFM
   generic map (
      DATA_WIDTH => FL_DATA_WIDTH,
      FL_BFM_ID => 00
   )
   port map (
      -- Common interface
      RESET           => reset,
      CLK             => clk,

      -- FrameLink input interface
      TX_DATA         => rx_data,
      TX_REM          => rx_rem,
      TX_SOF_N        => rx_sof_n,
      TX_EOF_N        => rx_eof_n,
      TX_SOP_N        => rx_sop_n,
      TX_EOP_N        => rx_eop_n,
      TX_SRC_RDY_N    => rx_src_rdy_n,
      TX_DST_RDY_N    => rx_dst_rdy_n
   ); 
   
	 -- -------------------------------------------------------------------------
   --                           Output FL_MONITOR
   -- -------------------------------------------------------------------------
   FL_MONITOR_I : entity work.MONITOR
   generic map (
      RX_TX_DATA_WIDTH => FL_DATA_WIDTH,
      FILE_NAME  => "./output/monitor",
      FRAME_PARTS => 1,
      RDY_DRIVER => RND
   )
   port map (
      -- Common interface
      FL_RESET        => reset,
      FL_CLK          => clk,

      -- FrameLink output interface
      RX_DATA         => tx_data,
      RX_REM          => tx_rem,
      RX_SOF_N        => tx_sof_n,
      RX_EOF_N        => tx_eof_n,
      RX_SOP_N        => tx_sop_n,
      RX_EOP_N        => tx_eop_n,
      RX_SRC_RDY_N    => tx_src_rdy_n,
      RX_DST_RDY_N    => tx_dst_rdy_n
   ); 
	 
   -- -------------------------------------------------------------------------
   --                           CLOCKs & RESETs
   -- -------------------------------------------------------------------------
   resetp : process
   begin
      reset <= '1', '0' after RESET_TIME;
      wait;
   end process;

   clk_genp: process
   begin
      clk  <= '1';
      wait for CLK_PERIOD/2;
      clk  <= '0';
      wait for CLK_PERIOD/2;
   end process;

   -- -----------------------------------------------------------------------
   --                             MI32 interface
   -- -----------------------------------------------------------------------

   mi32_dwr      <= (others => '0');
   mi32_addr     <= (others => '0');
   mi32_rd       <= '0';
   mi32_wr       <= '0';
   mi32_be       <= (others => '0');

   -- -----------------------------------------------------------------------
   --                                 Test
   -- -----------------------------------------------------------------------
   tb : process

   begin
      wait for RESET_TIME;

      report "========== start of core simulation ==========";
      SendWriteFile("./input/input_program_hex", RND, flCmd_0, 0);
      wait for 1200 us;
      --SendWriteFile("./input/input_program_hex", EVER, flCmd_0, 0);
      wait for 50us;--1200 us;
      --SendWriteFile("./input/input_program_hex", EVER, flCmd_0, 0);

      wait;

   end process;


end architecture;
